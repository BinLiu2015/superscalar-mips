��l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;    
 u s e   I E E E . N U M E R I C _ S T D _ U N S I G N E D . a l l ;  
  
 e n t i t y   a d d e r   i s   - -   a d d e r  
     p o r t ( a ,   b :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
               y :         o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   a d d e r   i s  
 b e g i n  
     y   < =   a   +   b ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;    
 u s e   I E E E . N U M E R I C _ S T D _ U N S I G N E D . a l l ;  
  
 e n t i t y   a l u   i s    
     p o r t ( a ,   b   :   i n   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         a l u c o n t r o l   :   i n           S T D _ L O G I C _ V E C T O R ( 2   d o w n t o   0 ) ;  
         r e s u l t           :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         z e r o               :   o u t         S T D _ L O G I C ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   a l u   i s  
     s i g n a l   c o n d i n v b ,   s u m   :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 b e g i n  
     c o n d i n v b   < =   n o t   b   w h e n   a l u c o n t r o l ( 2 )   e l s e   b ;  
     s u m             < =   a   +   c o n d i n v b   +   a l u c o n t r o l ( 2 ) ;  
      
     p r o c e s s ( a l l )   b e g i n  
         c a s e   a l u c o n t r o l ( 1   d o w n t o   0 )   i s  
             w h e n   " 0 0 "       = >   r e s u l t       < =   a   a n d   b ;    
             w h e n   " 0 1 "       = >   r e s u l t       < =   a   o r   b ;    
             w h e n   " 1 0 "       = >   r e s u l t       < =   s u m ;    
             w h e n   " 1 1 "       = >   r e s u l t       < =   ( 0   = >   s u m ( 3 1 ) ,   o t h e r s   = >   ' 0 ' ) ;    
             w h e n   o t h e r s   = >   r e s u l t   < =   ( o t h e r s   = >   ' X ' ) ;    
         e n d   c a s e ;  
     e n d   p r o c e s s ;  
      
     z e r o   < =   ' 1 '   w h e n   r e s u l t   =   X " 0 0 0 0 0 0 0 0 "   e l s e   ' 0 ' ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
  
 e n t i t y   a l u d e c   i s   - -   A L U   c o n t r o l   d e c o d e r  
     p o r t ( f u n c t   :   i n   S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
         a l u o p             :   i n     S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
         a l u c o n t r o l   :   o u t   S T D _ L O G I C _ V E C T O R ( 2   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   a l u d e c   i s  
 b e g i n  
     p r o c e s s ( a l l )   b e g i n  
         c a s e   a l u o p   i s  
                     w h e n   " 0 0 "           = >   a l u c o n t r o l   < =   " 0 1 0 " ;   - -   a d d   ( f o r   l w / s w / a d d i )  
                     w h e n   " 0 1 "           = >   a l u c o n t r o l   < =   " 1 1 0 " ;   - -   s u b   ( f o r   b e q )  
                     w h e n   " 1 1 "           = >   a l u c o n t r o l   < =   " 0 0 1 " ;   - -   o r   ( f o r   o r i )  
                     w h e n   o t h e r s       = >   c a s e   f u n c t   i s   - -   R - t y p e   i n s t r u c t i o n s  
                         w h e n   " 1 0 0 0 0 0 "   = >   a l u c o n t r o l   < =   " 0 1 0 " ;   - -   a d d    
                         w h e n   " 1 0 0 0 1 0 "   = >   a l u c o n t r o l   < =   " 1 1 0 " ;   - -   s u b  
                         w h e n   " 1 0 0 1 0 0 "   = >   a l u c o n t r o l   < =   " 0 0 0 " ;   - -   a n d  
                         w h e n   " 1 0 0 1 0 1 "   = >   a l u c o n t r o l   < =   " 0 0 1 " ;   - -   o r  
                         w h e n   " 1 0 1 0 1 0 "   = >   a l u c o n t r o l   < =   " 1 1 1 " ;   - -   s l t  
                         w h e n   o t h e r s       = >   a l u c o n t r o l       < =   " - - - " ;   - -   ? ? ?  
                 e n d   c a s e ;  
         e n d   c a s e ;  
     e n d   p r o c e s s ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
  
 e n t i t y   c o n t r o l l e r   i s   - -   s i n g l e   c y c l e   c o n t r o l   d e c o d e r  
 	 p o r t ( o p ,   f u n c t   :   i n   S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
 	 	 z e r o                               :   i n     S T D _ L O G I C ;  
 	 	 s t a l l 	 	 	       :   i n     S T D _ L O G I C ;  
 	 	 m e m t o r e g ,   m e m w r i t e   :   o u t   S T D _ L O G I C ;  
 	 	 p c s r c                             :   o u t   S T D _ L O G I C ;  
 	 	 a l u s r c                           :   o u t   S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 	 r e g d s t ,   r e g w r i t e       :   o u t   S T D _ L O G I C ;  
 	 	 j u m p                               :   o u t   S T D _ L O G I C ;  
 	 	 a l u c o n t r o l                   :   o u t   S T D _ L O G I C _ V E C T O R ( 2   d o w n t o   0 ) ) ;  
 e n d ;  
  
  
 a r c h i t e c t u r e   s t r u c t   o f   c o n t r o l l e r   i s  
 	 c o m p o n e n t   m a i n d e c  
 	 	 p o r t ( o p   :   i n   S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
 	 	 	 m e m t o r e g ,   m e m w r i t e   :   o u t   S T D _ L O G I C ;  
 	 	 	 b r a n c h                           :   o u t   S T D _ L O G I C ;  
 	 	 	 a l u s r c                           :   o u t   S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 	 	 r e g d s t ,   r e g w r i t e       :   o u t   S T D _ L O G I C ;  
 	 	 	 j u m p                               :   o u t   S T D _ L O G I C ;  
 	 	 	 a l u o p                             :   o u t   S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 	 	 b r a n c h N o t E q u a l           :   o u t   S T D _ L O G I C ) ;  
 	 e n d   c o m p o n e n t ;  
 	 c o m p o n e n t   a l u d e c  
 	 	 p o r t ( f u n c t   :   i n   S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
 	 	 	 a l u o p             :   i n     S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 	 	 a l u c o n t r o l   :   o u t   S T D _ L O G I C _ V E C T O R ( 2   d o w n t o   0 ) ) ;  
 	 e n d   c o m p o n e n t ;  
 	 s i g n a l   a l u o p                     :   S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 s i g n a l   b r a n c h                   :   S T D _ L O G I C ;  
 	 s i g n a l   b r a n c h N o t E q u a l   :   S T D _ L O G I C ;  
 	 s i g n a l   t m p _ m e m w r i t e   :   S T D _ L O G I C ;  
 	 s i g n a l   t m p _ r e g w r i t e   :   S T D _ L O G I C ;  
 b e g i n  
 	 	 m d   :   m a i n d e c   p o r t   m a p ( o p ,   m e m t o r e g ,   t m p _ m e m w r i t e ,   b r a n c h ,  
 	 	 	 a l u s r c ,   r e g d s t ,   t m p _ r e g w r i t e ,   j u m p ,   a l u o p ,   b r a n c h N o t E q u a l ) ;  
 	 	 a d   :   a l u d e c   p o r t   m a p ( f u n c t ,   a l u o p ,   a l u c o n t r o l ) ;  
 	  
 	 m e m w r i t e   < =   t m p _ m e m w r i t e   a n d   n o t   s t a l l ;  
 	 r e g w r i t e   < =   t m p _ r e g w r i t e   a n d   n o t   s t a l l ;  
 	 p c s r c   < =   ( b r a n c h   a n d   z e r o )   o r   ( b r a n c h N o t E q u a l   a n d   n o t   z e r o ) ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;   u s e   I E E E . S T D _ L O G I C _ A R I T H . a l l ;  
      
 e n t i t y   d a t a p a t h   i s   - -   M I P S   d a t a p a t h  
     p o r t ( c l k ,   r e s e t   :   i n   S T D _ L O G I C ;  
         m e m t o r e g ,   p c s r c       :   i n           S T D _ L O G I C ;  
         a l u s r c                         :   i n           S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
         r e g d s t                         :   i n           S T D _ L O G I C ;  
         j u m p                             :   i n           S T D _ L O G I C ;  
         a l u c o n t r o l                 :   i n           S T D _ L O G I C _ V E C T O R ( 2   d o w n t o   0 ) ;  
         z e r o                             :   o u t         S T D _ L O G I C ;  
         p c                                 :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         i n s t r                           :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         a l u o u t                         :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         w r i t e d a t a                   :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         r e a d d a t a                     :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         p c n e x t                         :   o u t         S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         w r i t e r e g                     :   o u t         S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
         r e s u l t                         :   o u t         S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         s r c a                             :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   s t r u c t   o f   d a t a p a t h   i s  
     c o m p o n e n t   a l u  
         p o r t ( a ,   b   :   i n   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
             a l u c o n t r o l   :   i n           S T D _ L O G I C _ V E C T O R ( 2   d o w n t o   0 ) ;  
             r e s u l t           :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
             z e r o               :   o u t         S T D _ L O G I C ) ;  
     e n d   c o m p o n e n t ;  
     - -   c o m p o n e n t   r e g f i l e  
     - -       p o r t ( c l k   :   i n   S T D _ L O G I C ;  
     - -           w e 3                       :   i n     S T D _ L O G I C ;  
     - -           r a 1 ,   r a 2 ,   w a 3   :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
     - -           w d 3                       :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
     - -           r d 1 ,   r d 2             :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
     - -   e n d   c o m p o n e n t ;  
     c o m p o n e n t   a d d e r  
         p o r t ( a ,   b   :   i n   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
             y   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
     e n d   c o m p o n e n t ;  
     c o m p o n e n t   s l 2  
         p o r t ( a   :   i n   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
             y   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
     e n d   c o m p o n e n t ;  
     c o m p o n e n t   s i g n e x t  
         p o r t ( a   :   i n   S T D _ L O G I C _ V E C T O R ( 1 5   d o w n t o   0 ) ;  
             y   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
     e n d   c o m p o n e n t ;  
     - -   c o m p o n e n t   f l o p r   g e n e r i c ( w i d t h   :         i n t e g e r ) ;  
     - -       p o r t ( c l k ,   r e s e t                               :   i n   S T D _ L O G I C ;  
     - -           d   :   i n     S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ;  
     - -           q   :   o u t   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ) ;  
     - -   e n d   c o m p o n e n t ;  
     c o m p o n e n t   m u x 2   g e n e r i c ( w i d t h   :         i n t e g e r ) ;  
         p o r t ( d 0 ,   d 1                                     :   i n   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ;  
             s   :   i n     S T D _ L O G I C ;  
             y   :   o u t   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ) ;  
     e n d   c o m p o n e n t ;    
     c o m p o n e n t   m u x 4   g e n e r i c   ( w i d t h   :         i n t e g e r ) ;  
         p o r t ( d 0 , d 1 , d 2 , d 3                             :   i n   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ;  
             s   :   i n     S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
             y   :   o u t   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ) ;  
     e n d   c o m p o n e n t ;  
     - -   s i g n a l   w r i t e r e g   :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
     s i g n a l   p c j u m p ,    
     p c n e x t b r ,   p c p l u s 4 ,    
     p c b r a n c h                                     :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
     s i g n a l   s i g n i m m ,   s i g n i m m s h   :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
     s i g n a l   s r c b                               :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 b e g i n  
     - -   n e x t   P C   l o g i c  
     p c j u m p   < =   p c p l u s 4 ( 3 1   d o w n t o   2 8 )   &   i n s t r ( 2 5   d o w n t o   0 )   &   " 0 0 " ;  
         - -   p c r e g       :   f l o p r   g e n e r i c   m a p ( 3 2 )   p o r t   m a p ( c l k ,   r e s e t ,   p c n e x t ,   p c ) ;    
         p c a d d 1     :   a d d e r   p o r t   m a p ( p c ,   X " 0 0 0 0 0 0 0 4 " ,   p c p l u s 4 ) ;  
         i m m s h       :   s l 2   p o r t   m a p ( s i g n i m m ,   s i g n i m m s h ) ;  
         p c a d d 2     :   a d d e r   p o r t   m a p ( p c p l u s 4 ,   s i g n i m m s h ,   p c b r a n c h ) ;  
         p c b r m u x   :   m u x 2   g e n e r i c   m a p ( 3 2 )   p o r t   m a p ( p c p l u s 4 ,   p c b r a n c h ,    
             p c s r c ,   p c n e x t b r ) ;  
         p c m u x   :   m u x 2   g e n e r i c   m a p ( 3 2 )   p o r t   m a p ( p c n e x t b r ,   p c j u m p ,   j u m p ,   p c n e x t ) ;  
      
     - -   r e g i s t e r   f i l e   l o g i c  
         - -   r f   :   r e g f i l e   p o r t   m a p ( c l k ,   r e g w r i t e ,   i n s t r ( 2 5   d o w n t o   2 1 ) ,    
         - -       i n s t r ( 2 0   d o w n t o   1 6 ) ,   w r i t e r e g ,   r e s u l t ,   s r c a ,    
         - -       w r i t e d a t a ) ;  
         w r m u x   :   m u x 2   g e n e r i c   m a p ( 5 )   p o r t   m a p ( i n s t r ( 2 0   d o w n t o   1 6 ) ,    
             i n s t r ( 1 5   d o w n t o   1 1 ) ,    
             r e g d s t ,   w r i t e r e g ) ;  
         r e s m u x   :   m u x 2   g e n e r i c   m a p ( 3 2 )   p o r t   m a p ( a l u o u t ,   r e a d d a t a ,    
             m e m t o r e g ,   r e s u l t ) ;  
         s e   :   s i g n e x t   p o r t   m a p ( i n s t r ( 1 5   d o w n t o   0 ) ,   s i g n i m m ) ;  
      
     - -   A L U   l o g i c  
         s r c b m u x   :   m u x 4   g e n e r i c   m a p ( 3 2 )  
         p o r t   m a p (  
             d 0   = >   w r i t e d a t a ,  
             d 1   = >   " 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 " ,  
             d 2   = >   s i g n i m m ,  
             d 3   = >   " 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 "   &   i n s t r ( 1 5   d o w n t o   0 ) ,  
             s     = >   a l u s r c ,  
             y     = >   s r c b  
         ) ;  
         m a i n a l u   :   a l u   p o r t   m a p ( s r c a ,   s r c b ,   a l u c o n t r o l ,   a l u o u t ,   z e r o ) ;  
 e n d ;  
 l i b r a r y   I E E E ;    
 u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;   u s e   S T D . T E X T I O . a l l ;  
 u s e   I E E E . N U M E R I C _ S T D _ U N S I G N E D . a l l ;    
  
 e n t i t y   d m e m   i s   - -   d a t a   m e m o r y  
 	 p o r t ( c l k 	   :   i n     S T D _ L O G I C ;  
 	 	   w e 1 	   :   i n     S T D _ L O G I C ;  
 	 	   a 1 	 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	   w d 1 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	   r d 1   	   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	   w e 2 	   :   i n     S T D _ L O G I C ;  
 	 	   a 2 	   	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	   w d 2 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	   r d 2     	   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	   w e 3 	   :   i n     S T D _ L O G I C ;  
 	 	   a 3 	 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	   w d 3 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	   r d 3   	   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   d m e m   i s  
  
 b e g i n  
 	 p r o c e s s   i s  
 	 	 t y p e   r a m t y p e   i s   a r r a y   ( 6 3   d o w n t o   0 )   o f   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 v a r i a b l e   m e m :   r a m t y p e ;  
 	 b e g i n  
 	 	 - -   r e a d   o r   w r i t e   m e m o r y  
 	 	 l o o p  
 	 	 	 i f   c l k ' e v e n t   a n d   c l k   =   ' 1 '   t h e n  
 	 	 	 	 i f   ( w e 1   =   ' 1 '   a n d   ( ( ( a 1   / =   a 2 )   o r   ( w e 2   =   ' 0 ' ) )   a n d   ( ( a 1   / =   a 3 )   o r   ( w e 3   =   ' 0 ' ) ) ) )   t h e n    
 	 	 	 	 	 m e m ( t o _ i n t e g e r ( a 1 ( 7   d o w n t o   2 ) ) )   : =   w d 1 ;  
 	 	 	 	 e n d   i f ;  
 	 	 	 	 i f   ( w e 2   =   ' 1 '   a n d   ( ( a 2   / =   a 3 )   o r   ( w e 3   =   ' 0 ' ) ) )   t h e n    
 	 	 	 	 	 m e m ( t o _ i n t e g e r ( a 2 ( 7   d o w n t o   2 ) ) )   : =   w d 2 ;  
 	 	 	 	 e n d   i f ;  
 	 	 	 	 i f   ( w e 3   =   ' 1 ' )   t h e n  
 	 	 	 	 	 m e m ( t o _ i n t e g e r ( a 3 ( 7   d o w n t o   2 ) ) )   : =   w d 3 ;  
 	 	 	 	 e n d   i f ;  
 	 	 	 e n d   i f ;  
 	 	 	 r d 1   < =   m e m ( t o _ i n t e g e r ( a 1 ( 7   d o w n t o   2 ) ) ) ;    
 	 	 	 r d 2   < =   m e m ( t o _ i n t e g e r ( a 2 ( 7   d o w n t o   2 ) ) ) ;    
 	 	 	 r d 3   < =   m e m ( t o _ i n t e g e r ( a 3 ( 7   d o w n t o   2 ) ) ) ;   	 	 	  
 	 	 	 w a i t   o n   c l k ,   a 1 ,   a 2 ,   a 3 ;  
 	 	 e n d   l o o p ;  
 	 	  
 	 e n d   p r o c e s s ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;     u s e   I E E E . S T D _ L O G I C _ A R I T H . a l l ;  
  
 e n t i t y   f l o p r   i s   - -   f l i p - f l o p   w i t h   s y n c h r o n o u s   r e s e t  
     g e n e r i c ( w i d t h :   i n t e g e r ) ;  
     p o r t ( c l k ,   r e s e t :   i n     S T D _ L O G I C ;  
               d :                     i n     S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ;  
               q :                     o u t   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   a s y n c h r o n o u s   o f   f l o p r   i s  
 b e g i n  
     p r o c e s s ( c l k ,   r e s e t )   b e g i n  
         i f   r e s e t   t h e n     q   < =   ( o t h e r s   = >   ' 0 ' ) ;  
         e l s i f   r i s i n g _ e d g e ( c l k )   t h e n  
             q   < =   d ;  
         e n d   i f ;  
     e n d   p r o c e s s ;  
 e n d ;  
 l i b r a r y   I E E E ;    
 u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;   u s e   I E E E . N U M E R I C _ S T D _ U N S I G N E D . a l l ;  
  
 e n t i t y   h a z a r d u n i t   i s    
 	 p o r t ( c l k ,   r e s e t :   i n   S T D _ L O G I C ;  
 	 	 	 p c                               :   o u t     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 p c 1                             :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 i n s t r 1                       :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 j u m p 1                         :   i n       S T D _ L O G I C ;  
 	 	 	 p c s r c 1                       :   i n       S T D _ L O G I C ;  
 	 	 	 w r i t e r e g 1                 :   i n       S T D _ L O G I C ;  
 	 	 	 p c a d d r 1                     :   o u t     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 p c 2                             :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 i n s t r 2                       :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 j u m p 2                         :   i n       S T D _ L O G I C ;  
 	 	 	 p c s r c 2                       :   i n       S T D _ L O G I C ;  
 	 	 	 w r i t e r e g 2                 :   i n       S T D _ L O G I C ;  
 	 	 	 p c a d d r 2                     :   o u t     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 s t a l l 2                       :   b u f f e r     S T D _ L O G I C ;  
 	 	 	 p c 3                             :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 i n s t r 3                       :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 j u m p 3                         :   i n       S T D _ L O G I C ;  
 	 	 	 p c s r c 3                       :   i n       S T D _ L O G I C ;  
 	 	 	 w r i t e r e g 3                 :   i n       S T D _ L O G I C ;  
 	 	 	 p c a d d r 3                     :   o u t     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 s t a l l 3                       :   o u t     S T D _ L O G I C ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   t e s t   o f   h a z a r d u n i t   i s  
 	 c o m p o n e n t   j u m p s t a l l e r  
 	 	 p o r t ( j u m p 1 ,   p c s r c 1 :   i n   S T D _ L O G I C ;  
 	 	 	 j u m p 2 ,   p c s r c 2 :   i n   S T D _ L O G I C ;  
 	 	 	 j u m p 3 ,   p c s r c 3 :   i n   S T D _ L O G I C ;  
 	 	 	 s t a l l 2 ,   s t a l l 3 :   o u t   S T D _ L O G I C ) ;  
 	 e n d   c o m p o n e n t ;  
 	 c o m p o n e n t   m e m o r y s t a l l e r  
                 p o r t ( o p 1         :   i n     S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
                         b a s e r e g 1     :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
                         o f f s e t 1       :   i n     S T D _ L O G I C _ V E C T O R ( 1 5   d o w n t o   0 ) ;  
                         o p 2               :   i n     S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
                         b a s e r e g 2     :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
                         o f f s e t 2       :   i n     S T D _ L O G I C _ V E C T O R ( 1 5   d o w n t o   0 ) ;  
                         o p 3               :   i n     S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
                         b a s e r e g 3     :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
                         o f f s e t 3       :   i n     S T D _ L O G I C _ V E C T O R ( 1 5   d o w n t o   0 ) ;  
                         s t a l l 2 ,   s t a l l 3 :   o u t   S T D _ L O G I C ) ;              
     	 e n d   c o m p o n e n t ;  
 	 c o m p o n e n t   r e g s t a l l e r  
                 p o r t ( w r i t e r e g 1         :   i n     S T D _ L O G I C ;      
                           i n s t r 1                 :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
                           w r i t e r e g 2           :   i n     S T D _ L O G I C ;  
                           i n s t r 2                 :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
                           w r i t e r e g 3           :   i n     S T D _ L O G I C ;  
                           i n s t r 3                 :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
                           s t a l l 2 ,   s t a l l 3 :   o u t   S T D _ L O G I C ) ;              
     	 e n d   c o m p o n e n t ;  
         c o m p o n e n t   f l o p r   g e n e r i c ( w i d t h   :         i n t e g e r ) ;  
 	 	 p o r t ( c l k ,   r e s e t                               :   i n   S T D _ L O G I C ;  
 	 	 d   :   i n     S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ;  
 	 	 q   :   o u t   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ) ;  
     	 e n d   c o m p o n e n t ;  
  
 	 s i g n a l   p c n e x t ,   i n s t r ,   r e a d d a t a ,   r e s u l t ,   s r c a :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
         s i g n a l   j u m p _ s t a l l 2 ,   m e m _ s t a l l 2 ,   r e g _ s t a l l 2 :   S T D _ L O G I C ;  
         s i g n a l   j u m p _ s t a l l 3 ,   m e m _ s t a l l 3 ,   r e g _ s t a l l 3 :   S T D _ L O G I C ;  
 b e g i n  
         s t a l l 2   < =   j u m p _ s t a l l 2   o r   m e m _ s t a l l 2   o r   r e g _ s t a l l 2 ;  
         s t a l l 3   < =   j u m p _ s t a l l 3   o r   m e m _ s t a l l 3   o r   r e g _ s t a l l 3   o r   s t a l l 2 ;  
  
         p c n e x t   < =   p c 1   w h e n   s t a l l 2   a n d   s t a l l 3   e l s e  
                             p c 2   w h e n   s t a l l 3   e l s e  
                             p c 3 ;  
  
         p c a d d r 1   < =   p c ;  
         p c a d d r 2   < =   p c   +   " 1 0 0 " ;  
         p c a d d r 3   < =   p c   +   " 1 0 0 0 " ;  
  
  
         j s :   j u m p s t a l l e r   p o r t   m a p (  
                 j u m p 1   = >   j u m p 1 ,  
                 p c s r c 1   = >   p c s r c 1 ,  
                 j u m p 2   = >   j u m p 2 ,  
                 p c s r c 2   = >   p c s r c 2 ,  
                 j u m p 3   = >   j u m p 3 ,  
                 p c s r c 3   = >   p c s r c 3 ,  
                 s t a l l 2   = >   j u m p _ s t a l l 2 ,  
                 s t a l l 3   = >   j u m p _ s t a l l 3  
                 ) ;  
  
         r s :   r e g s t a l l e r   p o r t   m a p (  
                 w r i t e r e g 1   = >   w r i t e r e g 1 ,  
                 i n s t r 1   = >   i n s t r 1 ,  
                 w r i t e r e g 2   = >   w r i t e r e g 2 ,  
                 i n s t r 2   = >   i n s t r 2 ,  
                 w r i t e r e g 3   = >   w r i t e r e g 3 ,  
                 i n s t r 3   = >   i n s t r 3 ,  
                 s t a l l 2   = >   r e g _ s t a l l 2 ,  
                 s t a l l 3   = >   r e g _ s t a l l 3  
                 ) ;  
          
         m s :   m e m o r y s t a l l e r   p o r t   m a p (  
                 o p 1   = >   i n s t r 1 ( 3 1   d o w n t o   2 6 ) ,  
                 b a s e r e g 1   = >   i n s t r 1 ( 2 5   d o w n t o   2 1 ) ,  
                 o f f s e t 1   = >   i n s t r 1 ( 1 5   d o w n t o   0 ) ,  
                 o p 2   = >   i n s t r 2 ( 3 1   d o w n t o   2 6 ) ,  
                 b a s e r e g 2   = >   i n s t r 2 ( 2 5   d o w n t o   2 1 ) ,  
                 o f f s e t 2   = >   i n s t r 2 ( 1 5   d o w n t o   0 ) ,  
                 o p 3   = >   i n s t r 3 ( 3 1   d o w n t o   2 6 ) ,  
                 b a s e r e g 3   = >   i n s t r 3 ( 2 5   d o w n t o   2 1 ) ,  
                 o f f s e t 3   = >   i n s t r 3 ( 1 5   d o w n t o   0 ) ,  
                 s t a l l 2   = >   m e m _ s t a l l 2 ,  
                 s t a l l 3   = >   m e m _ s t a l l 3  
         ) ;  
  
         p c r e g :   f l o p r   g e n e r i c   m a p ( 3 2 )   p o r t   m a p ( c l k ,   r e s e t ,   p c n e x t ,   p c ) ;    
 e n d ;  
 l i b r a r y   I E E E ;    
 u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;   u s e   S T D . T E X T I O . a l l ;  
 u s e   I E E E . N U M E R I C _ S T D _ U N S I G N E D . a l l ;    
  
 e n t i t y   i m e m   i s   - -   i n s t r u c t i o n   m e m o r y  
 	 p o r t ( a :   i n   S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
 	 	 r d 1 :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 r d 2 :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 r d 3 :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   i m e m   i s  
 b e g i n  
 	 p r o c e s s   i s  
 	 	 f i l e   m e m _ f i l e                           :   T E X T ;  
 	 	 v a r i a b l e   L                                 :   l i n e ;  
 	 	 v a r i a b l e   c h                               :   c h a r a c t e r ;  
 	 	 v a r i a b l e   i ,   i n d e x ,   r e s u l t   :   i n t e g e r ;  
 	 	 t y p e   r a m t y p e   i s   a r r a y   ( 6 3   d o w n t o   0 )   o f   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 v a r i a b l e   m e m :   r a m t y p e ;  
 	 b e g i n  
 	 	 - -   i n i t i a l i z e   m e m o r y   f r o m   f i l e  
 	 	 f o r   i   i n   0   t o   6 3   l o o p   - -   s e t   a l l   c o n t e n t s   l o w  
 	 	 	 m e m ( i )   : =   ( o t h e r s   = >   ' 0 ' ) ;  
 	 	 e n d   l o o p ;  
 	 	 i n d e x   : =   0 ;  
 	 	 F I L E _ O P E N ( m e m _ f i l e ,   " C : \ U s e r s \ a g o d i n h o \ D o c u m e n t s \ A r q u i t e t u r a 2 \ m e m f i l e 3 . d a t " ,   R E A D _ M O D E ) ;  
 	 	 w h i l e   n o t   e n d f i l e ( m e m _ f i l e )   l o o p  
 	 	 r e a d l i n e ( m e m _ f i l e ,   L ) ;  
 	 	 r e s u l t   : =   0 ;  
 	 	 f o r   i   i n   1   t o   8   l o o p  
 	 	 	 r e a d ( L ,   c h ) ;  
 	 	 	 i f   ' 0 '   < =   c h   a n d   c h   < =   ' 9 '   t h e n    
 	 	 	 	 r e s u l t   : =   c h a r a c t e r ' p o s ( c h )   -   c h a r a c t e r ' p o s ( ' 0 ' ) ;  
 	 	 	 e l s i f   ' a '   < =   c h   a n d   c h   < =   ' f '   t h e n  
 	 	 	 	 r e s u l t   : =   c h a r a c t e r ' p o s ( c h )   -   c h a r a c t e r ' p o s ( ' a ' ) + 1 0 ;  
 	 	 	 e l s e   r e p o r t   " F o r m a t   e r r o r   o n   l i n e   "   &   i n t e g e r ' i m a g e ( i n d e x )  
 	 	 	 	 s e v e r i t y   e r r o r ;  
 	 	 	 e n d   i f ;  
 	 	 	 m e m ( i n d e x ) ( 3 5 - i * 4   d o w n t o   3 2 - i * 4 )   : =   t o _ s t d _ l o g i c _ v e c t o r ( r e s u l t , 4 ) ;  
 	 	 e n d   l o o p ;  
 	 	 i n d e x   : =   i n d e x   +   1 ;  
 	 e n d   l o o p ;  
 	  
 	 - -   r e a d   m e m o r y  
 	 l o o p  
 	 	 r d 1   < =   m e m ( t o _ i n t e g e r ( a ) ) ;  
 	 	 r d 2   < =   m e m ( t o _ i n t e g e r ( a )   +   1 ) ;  
 	 	 r d 3   < =   m e m ( t o _ i n t e g e r ( a )   +   2 ) ;  
 	 	 w a i t   o n   a ;  
 	 e n d   l o o p ;  
 e n d   p r o c e s s ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
  
 e n t i t y   j u m p s t a l l e r   i s  
     p o r t ( j u m p 1 ,   p c s r c 1 :   i n   S T D _ L O G I C ;  
               j u m p 2 ,   p c s r c 2 :   i n   S T D _ L O G I C ;  
               j u m p 3 ,   p c s r c 3 :   i n   S T D _ L O G I C ;  
               s t a l l 2 ,   s t a l l 3 :   o u t   S T D _ L O G I C ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   j u m p s t a l l e r   i s  
 b e g i n  
     s t a l l 2   < =   j u m p 1   o r   p c s r c 1 ;    
     s t a l l 3   < =   j u m p 2   o r   p c s r c 2   o r   j u m p 1   o r   p c s r c 1 ;    
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
  
 e n t i t y   m a i n d e c   i s   - -   m a i n   c o n t r o l   d e c o d e r  
 	 p o r t ( o p   :   i n   S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
 	 	 m e m t o r e g ,   m e m w r i t e   :   o u t   S T D _ L O G I C ;  
 	 	 b r a n c h                           :   o u t   S T D _ L O G I C ;    
 	 	 a l u s r c                           :   o u t   S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 	 r e g d s t ,   r e g w r i t e       :   o u t   S T D _ L O G I C ;  
 	 	 j u m p                               :   o u t   S T D _ L O G I C ;  
 	 	 a l u o p                             :   o u t   S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 	 b r a n c h N o t E q u a l           :   o u t   S T D _ L O G I C ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   m a i n d e c   i s  
 	 s i g n a l   c o n t r o l s   :   S T D _ L O G I C _ V E C T O R ( 1 0   d o w n t o   0 ) ;  
 b e g i n  
 	 p r o c e s s ( a l l )   b e g i n  
 	 	 c a s e   o p   i s  
 	 	 	   w h e n   " 0 0 0 0 0 0 "   = >   c o n t r o l s   < =   " 1 1 0 0 0 0 0 0 1 0 0 " ;   - -   R T Y P E  
 	 	 	   w h e n   " 1 0 0 0 1 1 "   = >   c o n t r o l s   < =   " 1 0 1 0 0 0 1 0 0 0 0 " ;   - -   L W  
 	 	 	   w h e n   " 1 0 1 0 1 1 "   = >   c o n t r o l s   < =   " 0 0 1 0 0 1 0 0 0 0 0 " ;   - -   S W  
 	 	 	   w h e n   " 0 0 0 1 0 0 "   = >   c o n t r o l s   < =   " 0 0 0 0 1 0 0 0 0 1 0 " ;   - -   B E Q  
 	 	 	   w h e n   " 0 0 0 1 0 1 "   = >   c o n t r o l s   < =   " 0 0 0 0 1 0 0 0 0 1 1 " ;   - -   B N E  
 	 	 	   w h e n   " 0 0 1 0 0 0 "   = >   c o n t r o l s   < =   " 1 0 1 0 0 0 0 0 0 0 0 " ;   - -   A D D I  
 	 	 	   w h e n   " 0 0 0 0 1 0 "   = >   c o n t r o l s   < =   " 0 0 0 0 0 0 0 1 0 0 0 " ;   - -   J  
 	 	 	   w h e n   " 0 0 1 1 0 1 "   = >   c o n t r o l s   < =   " 1 0 1 1 0 0 0 0 1 1 0 " ;   - -   O R I  
 	 	 	   w h e n   o t h e r s       = >   c o n t r o l s       < =   " - - - - - - - - - - - " ;   - -   i l l e g a l   o p  
 	 	 e n d   c a s e ;  
 	 e n d   p r o c e s s ;  
 	  
 	 ( r e g w r i t e ,   r e g d s t ,   a l u s r c ,   b r a n c h ,   m e m w r i t e ,  
 	 	 m e m t o r e g ,   j u m p ,   a l u o p ( 1   d o w n t o   0 ) ,   b r a n c h N o t E q u a l )   < =   c o n t r o l s ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
  
 e n t i t y   m e m o r y s t a l l e r   i s  
   p o r t ( o p 1               :   i n     S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
             b a s e r e g 1     :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
             o f f s e t 1       :   i n     S T D _ L O G I C _ V E C T O R ( 1 5   d o w n t o   0 ) ;  
             o p 2               :   i n     S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
             b a s e r e g 2     :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
             o f f s e t 2       :   i n     S T D _ L O G I C _ V E C T O R ( 1 5   d o w n t o   0 ) ;  
             o p 3               :   i n     S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
             b a s e r e g 3     :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
             o f f s e t 3       :   i n     S T D _ L O G I C _ V E C T O R ( 1 5   d o w n t o   0 ) ;  
             s t a l l 2 ,   s t a l l 3 :   o u t   S T D _ L O G I C ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   m e m o r y s t a l l e r   i s  
 b e g i n  
     s t a l l 2   < =   ' 1 '   w h e n   ( o p 1   =   " 1 0 1 0 1 1 "   a n d   o p 2   =   " 1 0 0 0 1 1 "   a n d   b a s e r e g 1   =   b a s e r e g 2   a n d   o f f s e t 1   =   o f f s e t 2 )   e l s e   ' 0 ' ;  
 	 s t a l l 3   < =   ' 1 '   w h e n   ( o p 2   =   " 1 0 1 0 1 1 "   a n d   o p 3   =   " 1 0 0 0 1 1 "   a n d   b a s e r e g 2   =   b a s e r e g 3   a n d   o f f s e t 2   =   o f f s e t 3 )   o r  
                                           ( o p 1   =   " 1 0 1 0 1 1 "   a n d   o p 3   =   " 1 0 0 0 1 1 "   a n d   b a s e r e g 1   =   b a s e r e g 3   a n d   o f f s e t 1   =   o f f s e t 3 )   e l s e   ' 0 ' ;  
 e n d ;    
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
  
 e n t i t y   m i p s   i s   - -   s i n g l e   c y c l e   M I P S   p r o c e s s o r  
 	 p o r t ( c l k ,   r e s e t   :   i n   S T D _ L O G I C ;  
 	 	 p c                                 :   i n   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 i n s t r                           :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 s t a l l 	 	 	     :   i n   S T D _ L O G I C ;  
 	 	 m e m w r i t e                     :   o u t   S T D _ L O G I C ;  
 	 	 a l u o u t 	 	 	     :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 w r i t e d a t a 	 	     :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 r e a d d a t a                     :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 p c n e x t                         :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 r e g w r i t e                     :   o u t   S T D _ L O G I C ;  
 	 	 w r i t e r e g                     :   o u t   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	 	 r e s u l t 	                     :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 s r c a                             :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 j u m p                             :   b u f f e r     S T D _ L O G I C ;  
 	 	 p c s r c                           :   b u f f e r     S T D _ L O G I C ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   s t r u c t   o f   m i p s   i s  
 	 c o m p o n e n t   c o n t r o l l e r  
 	 	 p o r t ( o p ,   f u n c t   :   i n   S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
 	 	 	 z e r o                               :   i n     S T D _ L O G I C ;  
 	 	 	 s t a l l 	 	 	       :   i n     S T D _ L O G I C ;  
 	 	 	 m e m t o r e g ,   m e m w r i t e   :   o u t   S T D _ L O G I C ;  
 	 	 	 p c s r c                             :   o u t   S T D _ L O G I C ;  
 	 	 	 a l u s r c                           :   o u t   S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 	 	 r e g d s t ,   r e g w r i t e       :   o u t   S T D _ L O G I C ;  
 	 	 	 j u m p                               :   o u t   S T D _ L O G I C ;  
 	 	 	 a l u c o n t r o l                   :   o u t   S T D _ L O G I C _ V E C T O R ( 2   d o w n t o   0 ) ) ;  
 	 e n d   c o m p o n e n t ;  
 	 c o m p o n e n t   d a t a p a t h  
 	 	 p o r t ( c l k ,   r e s e t   :   i n   S T D _ L O G I C ;  
 	 	 	 m e m t o r e g ,   p c s r c       :   i n           S T D _ L O G I C ;  
 	 	 	 a l u s r c                         :   i n           S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 	 	 r e g d s t                         :   i n           S T D _ L O G I C ;  
 	 	 	 j u m p   	 	 	     :   i n           S T D _ L O G I C ;  
 	 	 	 a l u c o n t r o l                 :   i n           S T D _ L O G I C _ V E C T O R ( 2   d o w n t o   0 ) ;  
 	 	 	 z e r o                             :   o u t         S T D _ L O G I C ;  
 	 	 	 p c                                 :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 i n s t r                           :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 a l u o u t 	 	 	     :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 w r i t e d a t a 	 	     :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 r e a d d a t a                     :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 p c n e x t                         :   o u t         S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 w r i t e r e g                     :   o u t         S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	 	 	 r e s u l t 	                     :   o u t         S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 s r c a                             :   i n           S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
 	 e n d   c o m p o n e n t ;  
 	  
 	 s i g n a l   a l u s r c                                                                     :   S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
 	 s i g n a l   m e m t o r e g ,   r e g d s t   	 	 	 	       :   S T D _ L O G I C ;  
 	 s i g n a l   z e r o                                                                         :   S T D _ L O G I C ;  
 	 s i g n a l   a l u c o n t r o l                                                             :   S T D _ L O G I C _ V E C T O R ( 2   d o w n t o   0 ) ;  
 b e g i n  
 	 	 c o n t   :   c o n t r o l l e r   p o r t   m a p ( i n s t r ( 3 1   d o w n t o   2 6 ) ,   i n s t r ( 5   d o w n t o   0 ) ,  
 	 	 	 z e r o ,   s t a l l ,   m e m t o r e g ,   m e m w r i t e ,   p c s r c ,   a l u s r c ,  
 	 	 	 r e g d s t ,   r e g w r i t e ,   j u m p ,   a l u c o n t r o l ) ;  
 	 	 d p   :   d a t a p a t h   p o r t   m a p ( c l k ,   r e s e t ,   m e m t o r e g ,   p c s r c ,   a l u s r c ,   r e g d s t ,  
 	 	 	 j u m p ,   a l u c o n t r o l ,   z e r o ,   p c ,   i n s t r ,  
 	 	 	 a l u o u t ,   w r i t e d a t a ,   r e a d d a t a ,   p c n e x t ,   w r i t e r e g ,   r e s u l t ,   s r c a ) ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
  
 e n t i t y   m u x 2   i s   - -   t w o - i n p u t   m u l t i p l e x e r  
     g e n e r i c ( w i d t h :   i n t e g e r ) ;  
     p o r t ( d 0 ,   d 1 :   i n     S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ;  
               s :             i n     S T D _ L O G I C ;  
               y :             o u t   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   m u x 2   i s  
 b e g i n  
     y   < =   d 1   w h e n   s   e l s e   d 0 ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
          
 e n t i t y   m u x 4   i s   - -   f o u r - i n p u t   m u l t i p l e x e r  
         g e n e r i c ( w i d t h         :         i n t e g e r ) ;  
         p o r t ( d 0 , d 1 , d 2 , d 3   :   i n   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ;  
                 s   :   i n     S T D _ L O G I C _ V E C T O R ( 1   d o w n t o   0 ) ;  
                 y   :   o u t   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   m u x 4   i s  
 b e g i n  
         y   < =   d 0   w h e n   s = " 0 0 "   e l s e  
                 d 1           w h e n   s = " 0 1 "   e l s e  
                 d 2           w h e n   s = " 1 0 "   e l s e  
                 d 3 ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;    
 u s e   I E E E . N U M E R I C _ S T D _ U N S I G N E D . a l l ;  
  
 e n t i t y   r e g f i l e   i s   - -   t h r e e - p o r t   r e g i s t e r   f i l e  
     p o r t ( c l k   :   i n   S T D _ L O G I C ;  
 	 	 	   w r i t e E n 1           	       :   i n     S T D _ L O G I C ;  
 	 	 	   r a 1 A ,   r a 1 B ,   w a 1       :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	 	 	   w r i t e d a t a 1       	       :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   r e a d 1 A ,   r e a d 1 B         :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   w r i t e E n 2           	       :   i n     S T D _ L O G I C ;  
 	 	 	   r a 2 A ,   r a 2 B ,   w a 2       :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	 	 	   w r i t e d a t a 2       	       :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   r e a d 2 A ,   r e a d 2 B         :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   w r i t e E n 3           	       :   i n     S T D _ L O G I C ;  
 	 	 	   r a 3 A ,   r a 3 B ,   w a 3       :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	 	 	   w r i t e d a t a 3       	       :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   r e a d 3 A ,   r e a d 3 B         :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   r e g f i l e   i s  
     t y p e   r a m t y p e   i s   a r r a y   ( 3 1   d o w n t o   0 )   o f   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
     s i g n a l   m e m :   r a m t y p e ;  
 b e g i n  
     - -   t h r e e - p o r t e d   r e g i s t e r   f i l e  
     - -   r e a d   t w o   p o r t s   c o m b i n a t i o n a l l y  
     - -   w r i t e   t h i r d   p o r t   o n   r i s i n g   e d g e   o f   c l o c k  
     - -   r e g i s t e r   0   h a r d w i r e d   t o   0  
     - -   n o t e :   f o r   p i p e l i n e d   p r o c e s s o r ,   w r i t e   t h i r d   p o r t  
     - -   o n   f a l l i n g   e d g e   o f   c l k  
     p r o c e s s ( c l k )   b e g i n  
         i f   r i s i n g _ e d g e ( c l k )   t h e n  
               i f   c l k ' e v e n t   a n d   c l k   =   ' 1 '   t h e n  
 	 	 	 	 i f   ( w r i t e E n 1   =   ' 1 '   a n d   ( ( ( w a 1   / =   w a 2 )   o r   ( w r i t e E n 2   =   ' 0 ' ) )   a n d   ( ( w a 1   / =   w a 3 )   o r   ( w r i t e E n 3   =   ' 0 ' ) ) ) )   t h e n    
 	 	 	 	 	 m e m ( t o _ i n t e g e r ( w a 1 ) )   < =   w r i t e d a t a 1 ;  
 	 	 	 	 e n d   i f ;  
 	 	 	 	 i f   ( w r i t e E n 2   =   ' 1 '   a n d   ( ( w a 2   / =   w a 3 )   o r   ( w r i t e E n 3   =   ' 0 ' ) ) )   t h e n    
 	 	 	 	 	 m e m ( t o _ i n t e g e r ( w a 2 ) )   < =   w r i t e d a t a 2 ;  
 	 	 	 	 e n d   i f ;  
 	 	 	 	 i f   ( w r i t e E n 3   =   ' 1 ' )   t h e n  
 	 	 	 	 	 m e m ( t o _ i n t e g e r ( w a 3 ) )   < =   w r i t e d a t a 3 ;  
 	 	 	 	 e n d   i f ;  
 	 	 	 e n d   i f ;  
         e n d   i f ;  
     e n d   p r o c e s s ;  
     p r o c e s s ( a l l )   b e g i n  
         i f   ( t o _ i n t e g e r ( r a 1 A )   =   0 )   t h e n   r e a d 1 A   < =   X " 0 0 0 0 0 0 0 0 " ;   - -   r e g i s t e r   0   h o l d s   0  
         e l s e   r e a d 1 A   < =   m e m ( t o _ i n t e g e r ( r a 1 A ) ) ;  
         e n d   i f ;  
         i f   ( t o _ i n t e g e r ( r a 1 B )   =   0 )   t h e n   r e a d 1 B   < =   X " 0 0 0 0 0 0 0 0 " ;    
         e l s e   r e a d 1 B   < =   m e m ( t o _ i n t e g e r ( r a 1 B ) ) ;  
         e n d   i f ;  
  
         i f   ( t o _ i n t e g e r ( r a 2 A )   =   0 )   t h e n   r e a d 2 A   < =   X " 0 0 0 0 0 0 0 0 " ;   - -   r e g i s t e r   0   h o l d s   0  
         e l s e   r e a d 2 A   < =   m e m ( t o _ i n t e g e r ( r a 2 A ) ) ;  
         e n d   i f ;  
         i f   ( t o _ i n t e g e r ( r a 2 B )   =   0 )   t h e n   r e a d 2 B   < =   X " 0 0 0 0 0 0 0 0 " ;    
         e l s e   r e a d 2 B   < =   m e m ( t o _ i n t e g e r ( r a 2 B ) ) ;  
         e n d   i f ;  
  
         i f   ( t o _ i n t e g e r ( r a 3 A )   =   0 )   t h e n   r e a d 3 A   < =   X " 0 0 0 0 0 0 0 0 " ;   - -   r e g i s t e r   0   h o l d s   0  
         e l s e   r e a d 3 A   < =   m e m ( t o _ i n t e g e r ( r a 3 A ) ) ;  
         e n d   i f ;  
         i f   ( t o _ i n t e g e r ( r a 3 B )   =   0 )   t h e n   r e a d 3 B   < =   X " 0 0 0 0 0 0 0 0 " ;    
         e l s e   r e a d 3 B   < =   m e m ( t o _ i n t e g e r ( r a 3 B ) ) ;  
         e n d   i f ;  
          
     e n d   p r o c e s s ;  
 e n d ;  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
 u s e   I E E E . N U M E R I C _ S T D _ U N S I G N E D . a l l ;  
  
 e n t i t y   r e g s t a l l e r   i s  
     p o r t ( w r i t e r e g 1           :   i n     S T D _ L O G I C ;  
               i n s t r 1                 :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
               w r i t e r e g 2           :   i n     S T D _ L O G I C ;  
               i n s t r 2                 :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
               w r i t e r e g 3           :   i n     S T D _ L O G I C ;  
               i n s t r 3                 :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
               s t a l l 2 ,   s t a l l 3 :   o u t   S T D _ L O G I C ) ;    
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   r e g s t a l l e r   i s  
         s i g n a l   d e s t 1 :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
         s i g n a l   s r c A 2 :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
         s i g n a l   s r c B 2 :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
         s i g n a l   d e s t 2 :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
         s i g n a l   s r c A 3 :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
         s i g n a l   s r c B 3 :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 b e g i n  
  
         d e s t 1   < =   i n s t r 1 ( 1 5   d o w n t o   1 1 )   w h e n   i n s t r 1 ( 3 1   d o w n t o   2 6 )   =   " 0 0 0 0 0 0 "   e l s e   i n s t r 1 ( 2 0   d o w n t o   1 6 ) ;  
         s r c A 2   < =   i n s t r 2 ( 2 5   d o w n t o   2 1 ) ;  
         s r c B 2   < =   i n s t r 2 ( 2 0   d o w n t o   1 6 )   w h e n   i n s t r 2 ( 3 1   d o w n t o   2 6 )   =   " 0 0 0 0 0 0 "   e l s e   i n s t r 2 ( 2 5   d o w n t o   2 1 ) ;  
  
         d e s t 2   < =   i n s t r 2 ( 1 5   d o w n t o   1 1 )   w h e n   i n s t r 2 ( 3 1   d o w n t o   2 6 )   =   " 0 0 0 0 0 0 "   e l s e   i n s t r 2 ( 2 0   d o w n t o   1 6 ) ;  
         s r c A 3   < =   i n s t r 3 ( 2 5   d o w n t o   2 1 ) ;  
         s r c B 3   < =   i n s t r 3 ( 2 0   d o w n t o   1 6 )   w h e n   i n s t r 3 ( 3 1   d o w n t o   2 6 )   =   " 0 0 0 0 0 0 "   e l s e   i n s t r 3 ( 2 5   d o w n t o   2 1 ) ;  
  
         s t a l l 2   < =   ' 1 '   w h e n   ( w r i t e r e g 1   =   ' 1 '   a n d   ( d e s t 1   =   s r c A 2   o r   d e s t 1   =   s r c B 2 ) )   e l s e   ' 0 ' ;  
 s t a l l 3   < =   ' 1 '   w h e n   ( w r i t e r e g 2   =   ' 1 '   a n d   ( d e s t 2   =   s r c A 3   o r   d e s t 2   =   s r c B 3 ) )   o r  
                                               ( w r i t e r e g 1   =   ' 1 '   a n d   ( d e s t 1   =   s r c A 3   o r   d e s t 1   =   s r c B 3 ) )   e l s e   ' 0 ' ;  
 e n d ;  
  
 l i b r a r y   I E E E ;  
 u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
  
 e n t i t y   s i g n e x t   i s   - -   s i g n   e x t e n d e r  
     p o r t (  
         a :   i n     S T D _ L O G I C _ V E C T O R ( 1 5   d o w n t o   0 ) ;  
         y :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 )  
     ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   s i g n e x t   o f   s i g n e x t   i s  
 b e g i n  
     y   < =   " 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 "   &   a   w h e n   a ( 1 5 )   =   ' 1 '   e l s e   " 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 "   &   a ;    
 e n d ;  
  
 l i b r a r y   I E E E ;   u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;  
  
 e n t i t y   s l 2   i s   - -   s h i f t   l e f t   b y   2  
     p o r t ( a :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
               y :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   b e h a v e   o f   s l 2   i s  
 b e g i n  
     y   < =   a ( 2 9   d o w n t o   0 )   &   " 0 0 " ;  
 e n d ;  
 - -   m i p s . v h d  
 - -   F r o m   S e c t i o n   7 . 6   o f   D i g i t a l   D e s i g n   &   C o m p u t e r   A r c h i t e c t u r e  
 - -   U p d a t e d   t o   V H D L   2 0 0 8   2 6   J u l y   2 0 1 1   D a v i d _ H a r r i s @ h m c . e d u  
  
 l i b r a r y   I E E E ;    
 u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;   u s e   I E E E . N U M E R I C _ S T D _ U N S I G N E D . a l l ;  
  
 e n t i t y   t e s t b e n c h   i s  
 e n d ;  
  
 a r c h i t e c t u r e   t e s t   o f   t e s t b e n c h   i s  
     c o m p o n e n t   t o p  
         p o r t ( c l k ,   r e s e t   :   i n   S T D _ L O G I C ;    
             w r i t e d a t a 1 ,   d a t a a d r 1   :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
             w r i t e d a t a 2 ,   d a t a a d r 2   :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
             w r i t e d a t a 3 ,   d a t a a d r 3   :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
             m e m w r i t e 1                         :   b u f f e r   S T D _ L O G I C ;  
             m e m w r i t e 2                         :   b u f f e r   S T D _ L O G I C ;  
             m e m w r i t e 3                         :   b u f f e r   S T D _ L O G I C ) ;  
     e n d   c o m p o n e n t ;  
     s i g n a l   w r i t e d a t a 1 ,   d a t a a d r 1                                                 :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
     s i g n a l   w r i t e d a t a 2 ,   d a t a a d r 2                                                 :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
     s i g n a l   w r i t e d a t a 3 ,   d a t a a d r 3                                                 :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
     s i g n a l   c l k ,   r e s e t ,   m e m w r i t e 1 ,   m e m w r i t e 2 ,   m e m w r i t e 3   :   S T D _ L O G I C ;  
 b e g i n  
      
     - -   i n s t a n t i a t e   d e v i c e   t o   b e   t e s t e d  
         d u t   :   t o p   p o r t   m a p ( c l k ,   r e s e t ,    
             w r i t e d a t a 1 ,   d a t a a d r 1 ,  
             w r i t e d a t a 2 ,   d a t a a d r 2 ,  
             w r i t e d a t a 3 ,   d a t a a d r 3 ,  
             m e m w r i t e 1 ,  
             m e m w r i t e 2 ,  
             m e m w r i t e 3 ) ;  
      
     - -   G e n e r a t e   c l o c k   w i t h   1 0   n s   p e r i o d  
     p r o c e s s   b e g i n  
         c l k   < =   ' 1 ' ;  
         w a i t   f o r   5   n s ;    
         c l k   < =   ' 0 ' ;  
         w a i t   f o r   5   n s ;  
     e n d   p r o c e s s ;  
      
     - -   G e n e r a t e   r e s e t   f o r   f i r s t   t w o   c l o c k   c y c l e s  
     p r o c e s s   b e g i n  
         r e s e t   < =   ' 1 ' ;  
         w a i t   f o r   2 2   n s ;  
         r e s e t   < =   ' 0 ' ;  
         w a i t ;  
     e n d   p r o c e s s ;  
      
     - -   c h e c k   t h a t   - 3 3 0 2 2   g e t s   w r i t t e n   t o   a d d r e s s   8 4   a t   e n d   o f   p r o g r a m  
     p r o c e s s   ( c l k )   b e g i n  
         i f   ( c l k ' e v e n t   a n d   c l k   =   ' 0 '   a n d   m e m w r i t e 1   =   ' 1 ' )   t h e n  
             i f   ( t o _ i n t e g e r ( d a t a a d r 1 )   =   8 4   a n d   t o _ i n t e g e r ( w r i t e d a t a 1 )   =   - 3 3 0 2 2 )   t h e n    
                 r e p o r t   " N O   E R R O R S   :   S i m u l a t i o n   s u c c e e d e d 1 "   s e v e r i t y   f a i l u r e ;  
             e l s i f   ( d a t a a d r 1   / =   8 0 )   t h e n    
                 r e p o r t   " S i m u l a t i o n   f a i l e d "   s e v e r i t y   f a i l u r e ;  
             e n d   i f ;  
         e n d   i f ;  
          
         i f   ( c l k ' e v e n t   a n d   c l k   =   ' 0 '   a n d   m e m w r i t e 2   =   ' 1 ' )   t h e n  
             i f   ( t o _ i n t e g e r ( d a t a a d r 2 )   =   8 4   a n d   t o _ i n t e g e r ( w r i t e d a t a 2 )   =   - 3 3 0 2 2 )   t h e n    
                 r e p o r t   " N O   E R R O R S   :   S i m u l a t i o n   s u c c e e d e d 2 "   s e v e r i t y   f a i l u r e ;  
             e l s i f   ( d a t a a d r 2   / =   8 0 )   t h e n    
                 r e p o r t   " S i m u l a t i o n   f a i l e d "   s e v e r i t y   f a i l u r e ;  
             e n d   i f ;  
         e n d   i f ;  
          
         i f   ( c l k ' e v e n t   a n d   c l k   =   ' 0 '   a n d   m e m w r i t e 3   =   ' 1 ' )   t h e n  
             i f   ( t o _ i n t e g e r ( d a t a a d r 3 )   =   8 4   a n d   t o _ i n t e g e r ( w r i t e d a t a 3 )   =   - 3 3 0 2 2 )   t h e n    
                 r e p o r t   " N O   E R R O R S   :   S i m u l a t i o n   s u c c e e d e d 3 "   s e v e r i t y   f a i l u r e ;  
             e l s i f   ( d a t a a d r 3   / =   8 0 )   t h e n    
                 r e p o r t   " S i m u l a t i o n   f a i l e d "   s e v e r i t y   f a i l u r e ;  
             e n d   i f ;  
         e n d   i f ;  
     e n d   p r o c e s s ;  
 e n d ;  
 l i b r a r y   I E E E ;    
 u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . a l l ;   u s e   I E E E . N U M E R I C _ S T D _ U N S I G N E D . a l l ;  
  
 e n t i t y   t o p   i s   - -   t o p - l e v e l   d e s i g n   f o r   t e s t i n g  
 	 p o r t ( c l k ,   r e s e t :   i n   S T D _ L O G I C ;  
 	 	 w r i t e d a t a 1 ,   d a t a a d r 1 :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 w r i t e d a t a 2 ,   d a t a a d r 2 :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 w r i t e d a t a 3 ,   d a t a a d r 3 :   b u f f e r   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 m e m w r i t e 1                     :   b u f f e r   S T D _ L O G I C ;  
 	 	 m e m w r i t e 2                     :   b u f f e r   S T D _ L O G I C ;  
 	 	 m e m w r i t e 3                     :   b u f f e r   S T D _ L O G I C ) ;  
 e n d ;  
  
 a r c h i t e c t u r e   t e s t   o f   t o p   i s  
 	 c o m p o n e n t   m i p s    
 	 	 p o r t ( c l k ,   r e s e t :   i n   S T D _ L O G I C ;  
 	 	 	 p c                               :   i n   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 i n s t r                         :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 s t a l l 	 	 	   :   i n     S T D _ L O G I C ; 	 	 	  
 	 	 	 m e m w r i t e                   :   o u t   S T D _ L O G I C ;  
 	 	 	 a l u o u t 	 	 	   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 w r i t e d a t a 	 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 r e a d d a t a                   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 p c n e x t                       :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 r e g w r i t e                   :   o u t   S T D _ L O G I C ;  
 	 	 	 w r i t e r e g                   :   o u t   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	 	 	 r e s u l t 	                   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 s r c a                           :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 j u m p                           :   b u f f e r     S T D _ L O G I C ;  
 	 	 	 p c s r c                         :   b u f f e r     S T D _ L O G I C ) ;  
 	 e n d   c o m p o n e n t ;  
 	 c o m p o n e n t   h a z a r d u n i t    
 	 	 p o r t ( c l k ,   r e s e t :   i n   S T D _ L O G I C ;  
 	 	 	 p c                               :   o u t     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 p c 1                             :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 i n s t r 1                       :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 j u m p 1                         :   i n       S T D _ L O G I C ;  
 	 	 	 p c s r c 1                       :   i n       S T D _ L O G I C ;  
 	 	 	 w r i t e r e g 1                 :   i n       S T D _ L O G I C ;  
 	 	 	 p c a d d r 1                     :   o u t     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 p c 2                             :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 i n s t r 2                       :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 j u m p 2                         :   i n       S T D _ L O G I C ;  
 	 	 	 p c s r c 2                       :   i n       S T D _ L O G I C ;  
 	 	 	 w r i t e r e g 2                 :   i n       S T D _ L O G I C ;  
 	 	 	 p c a d d r 2                     :   o u t     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 s t a l l 2                       :   b u f f e r     S T D _ L O G I C ;  
 	 	 	 p c 3                             :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 i n s t r 3                       :   i n       S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 j u m p 3                         :   i n       S T D _ L O G I C ;  
 	 	 	 p c s r c 3                       :   i n       S T D _ L O G I C ;  
 	 	 	 w r i t e r e g 3                 :   i n       S T D _ L O G I C ;  
 	 	 	 p c a d d r 3                     :   o u t     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 s t a l l 3                       :   o u t     S T D _ L O G I C ) ;  
 	 e n d   c o m p o n e n t ;  
 	 c o m p o n e n t   f l o p r   g e n e r i c ( w i d t h   :         i n t e g e r ) ;  
 	 	 p o r t ( c l k ,   r e s e t                               :   i n   S T D _ L O G I C ;  
 	 	 d   :   i n     S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ;  
 	 	 q   :   o u t   S T D _ L O G I C _ V E C T O R ( w i d t h - 1   d o w n t o   0 ) ) ;  
     	 e n d   c o m p o n e n t ;  
 	 c o m p o n e n t   i m e m  
 	 	 p o r t ( a :   i n   S T D _ L O G I C _ V E C T O R ( 5   d o w n t o   0 ) ;  
 	 	 	 r d 1 :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 r d 2 :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	 r d 3 :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
 	 e n d   c o m p o n e n t ;  
 	 c o m p o n e n t   d m e m  
 	 	 p o r t ( c l k 	   :   i n     S T D _ L O G I C ;    
 	 	 	   w e 1 	   :   i n     S T D _ L O G I C ;  
 	 	 	   a 1 	 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   w d 1 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   r d 1   	   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   w e 2 	   :   i n     S T D _ L O G I C ;  
 	 	 	   a 2 	   	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   w d 2 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   r d 2     	   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   w e 3 	   :   i n     S T D _ L O G I C ;  
 	 	 	   a 3 	 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   w d 3 	   :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   r d 3   	   :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;  
 	 e n d   c o m p o n e n t ;  
 	 c o m p o n e n t   r e g f i l e  
 	 	 p o r t ( c l k   :   i n   S T D _ L O G I C ;  
 	 	 	   w r i t e E n 1           	       :   i n     S T D _ L O G I C ;  
 	 	 	   r a 1 A ,   r a 1 B ,   w a 1       :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	 	 	   w r i t e d a t a 1       	       :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   r e a d 1 A ,   r e a d 1 B         :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   w r i t e E n 2           	       :   i n     S T D _ L O G I C ;  
 	 	 	   r a 2 A ,   r a 2 B ,   w a 2       :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	 	 	   w r i t e d a t a 2       	       :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   r e a d 2 A ,   r e a d 2 B         :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   w r i t e E n 3           	       :   i n     S T D _ L O G I C ;  
 	 	 	   r a 3 A ,   r a 3 B ,   w a 3       :   i n     S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	 	 	   w r i t e d a t a 3       	       :   i n     S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 	 	   r e a d 3 A ,   r e a d 3 B         :   o u t   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ) ;      
     	 e n d   c o m p o n e n t ;  
 	 s i g n a l   p c :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
  
 	 s i g n a l   r e g w r i t e 1 ,   p c s r c 1 ,   j u m p 1 :   S T D _ L O G I C ;  
 	 s i g n a l   i n s t r 1 ,   p c a d d r 1 ,   r e a d d a t a 1 ,   p c 1 ,   r e s u l t 1 ,   s r c a 1 :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 s i g n a l   w r i t e r e g 1 :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 	  
 	 s i g n a l   r e g w r i t e 2 ,   p c s r c 2 ,   j u m p 2 ,   s t a l l 2 :   S T D _ L O G I C ;  
 	 s i g n a l   i n s t r 2 ,   p c a d d r 2 ,   r e a d d a t a 2 ,   p c 2 ,   r e s u l t 2 ,   s r c a 2 :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 s i g n a l   w r i t e r e g 2 :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
  
 	 s i g n a l   r e g w r i t e 3 ,   p c s r c 3 ,   j u m p 3 ,   s t a l l 3 :   S T D _ L O G I C ;  
 	 s i g n a l   i n s t r 3 ,   p c a d d r 3 ,   r e a d d a t a 3 ,   p c 3 ,   r e s u l t 3 ,   s r c a 3 :   S T D _ L O G I C _ V E C T O R ( 3 1   d o w n t o   0 ) ;  
 	 s i g n a l   w r i t e r e g 3 :   S T D _ L O G I C _ V E C T O R ( 4   d o w n t o   0 ) ;  
 b e g i n  
 	 - -   i n s t a n t i a t e   p r o c e s s o r   a n d   m e m o r i e s  
 	 m i p s 1 :   m i p s   p o r t   m a p ( c l k ,   r e s e t ,   p c a d d r 1 ,   i n s t r 1 ,   ' 0 ' ,   m e m w r i t e 1 ,   d a t a a d r 1 ,  
 	 	 w r i t e d a t a 1 ,   r e a d d a t a 1 ,   p c 1 ,   r e g w r i t e 1 ,   w r i t e r e g 1 ,   r e s u l t 1 ,   s r c a 1 ,   j u m p 1 ,   p c s r c 1 ) ;  
 	  
 	 m i p s 2 :   m i p s   p o r t   m a p ( c l k ,   r e s e t ,   p c a d d r 2 ,   i n s t r 2 ,   s t a l l 2 ,   m e m w r i t e 2 ,   d a t a a d r 2 ,  
 	 	 w r i t e d a t a 2 ,   r e a d d a t a 2 ,   p c 2 ,   r e g w r i t e 2 ,   w r i t e r e g 2 ,   r e s u l t 2 ,   s r c a 2 ,   j u m p 2 ,   p c s r c 2 ) ;  
 	  
 	 m i p s 3 :   m i p s   p o r t   m a p ( c l k ,   r e s e t ,   p c a d d r 3 ,   i n s t r 3 ,   s t a l l 3 ,   m e m w r i t e 3 ,   d a t a a d r 3 ,  
 	 	 w r i t e d a t a 3 ,   r e a d d a t a 3 ,   p c 3 ,   r e g w r i t e 3 ,   w r i t e r e g 3 ,   r e s u l t 3 ,   s r c a 3 ,   j u m p 3 ,   p c s r c 3 ) ;  
  
 	  
 	 i m e m 1 :   i m e m   p o r t   m a p ( p c ( 7   d o w n t o   2 ) ,   i n s t r 1 ,   i n s t r 2 ,   i n s t r 3 ) ;  
  
 	 d m e m 1 :   d m e m   p o r t   m a p ( c l k ,   m e m w r i t e 1 ,   d a t a a d r 1 ,   w r i t e d a t a 1 ,   r e a d d a t a 1 ,  
 	 	 	 	 	 	 	     m e m w r i t e 2 ,   d a t a a d r 2 ,   w r i t e d a t a 2 ,   r e a d d a t a 2 ,  
 	 	 	 	 	 	 	     m e m w r i t e 3 ,   d a t a a d r 3 ,   w r i t e d a t a 3 ,   r e a d d a t a 3 ) ;  
 	  
  
 	 r f :   r e g f i l e   p o r t   m a p ( c l k ,    
 	 	 r e g w r i t e 1 ,   i n s t r 1 ( 2 5   d o w n t o   2 1 ) ,   i n s t r 1 ( 2 0   d o w n t o   1 6 ) ,   w r i t e r e g 1 ,   r e s u l t 1 ,   s r c a 1 ,   w r i t e d a t a 1 ,  
 	 	 r e g w r i t e 2 ,   i n s t r 2 ( 2 5   d o w n t o   2 1 ) ,   i n s t r 2 ( 2 0   d o w n t o   1 6 ) ,   w r i t e r e g 2 ,   r e s u l t 2 ,   s r c a 2 ,   w r i t e d a t a 2 ,  
 	 	 r e g w r i t e 3 ,   i n s t r 3 ( 2 5   d o w n t o   2 1 ) ,   i n s t r 3 ( 2 0   d o w n t o   1 6 ) ,   w r i t e r e g 3 ,   r e s u l t 3 ,   s r c a 3 ,   w r i t e d a t a 3 ) ;  
  
 	 h a z a r d :   h a z a r d u n i t   p o r t   m a p (  
 	 	 c l k ,   r e s e t ,   p c ,    
 	 	 p c 1 ,   i n s t r 1 ,   j u m p 1 ,   p c s r c 1 ,   r e g w r i t e 1 ,   p c a d d r 1 ,    
 	 	 p c 2 ,   i n s t r 2 ,   j u m p 2 ,   p c s r c 2 ,   r e g w r i t e 2 ,   p c a d d r 2 ,   s t a l l 2 ,    
 	 	 p c 3 ,   i n s t r 3 ,   j u m p 3 ,   p c s r c 3 ,   r e g w r i t e 3 ,   p c a d d r 3 ,   s t a l l 3 ) ;  
  
 e n d ;  
 